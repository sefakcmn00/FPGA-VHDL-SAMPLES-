
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity KOD is
    Port ( CLK : in  STD_LOGIC_VECTOR (1 downto 0)
	        basla: in std_logic;
	  );
end KOD;

architecture Behavioral of KOD is
signal count:integer 
begin


end Behavioral;

